library IEEE;
use IEEE.std_logic_1164.all;

entity hw01-1 is
    port(A,B,C,D : in std_logic;
        Z : out std_logic);
end hw01-1;

architecture structure of hw01-1 is
signal 